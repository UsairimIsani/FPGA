--www.21eda.net
--Email: sz21eda@126.com
--NET "key_data<0>"  LOC = "P111"  ;  K1
--NET "key_data<1>"  LOC = "P112"  ;  K2
--NET "key_data<2>"  LOC = "P114"  ;  K3
--NET "key_data<3>"  LOC = "P15"  ;   K4
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity KEY_LED is
PORT ( key_data  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);     --KEY input
       LED7      : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);     --
       LED7S     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)  ) ; --Digital tube display
end KEY_LED;

architecture Behavioral of KEY_LED is
 signal led_temp: std_logic_vector(3 downto 0);
 BEGIN 
  PROCESS( key_data ) 
  BEGIN 
     LED7 <="00000000" ;
     led_temp<= key_data ;
  CASE  led_temp  IS 
   WHEN "1110" =>  LED7S <= "11111001";    --  1
   WHEN "1101" =>  LED7S <= "10100100";    --  2
   WHEN "1011" =>  LED7S <= "10110000";    --  3
   WHEN "0111" =>  LED7S <= "10011001";    --  4
   WHEN OTHERS =>  LED7S <= "10000000";    --  8  --not key input display 8
   END CASE ; 
  END PROCESS ; 
  
end Behavioral;
