--www.21eda.net
--Email: sz21eda@126.com
-- VGA display 21EDA����
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LCD_VGA is

Port (     clk50_in : in std_logic;      --clk50M
           Red_out : out std_logic;      --R 
           Green_out : out std_logic;    --G
           Blue_out : out std_logic;     --B
           hs_out : out std_logic;       --hs clk
           vs_out : out std_logic);      --vs clk
end LCD_VGA;

architecture Behavioral of LCD_VGA is
signal Clk25					: std_logic; 
		signal Horizontal_Counter	: std_logic_vector (9 downto 0); 
		signal Vertical_Counter		: std_logic_vector (9 downto 0); 
 
begin 
--Generate 25Mhz Clock 
process (clk50_in) 
begin 
	if clk50_in'event and clk50_in='1' then 
	  if (Clk25 = '0')then 
	    Clk25 <= '1' after 2 ns; 
	  else 
	    Clk25 <= '0' after 2 ns; 
		end if; 
	end if; 
end process;		   
 
process (Clk25) 
TYPE Screen_Line1 is ARRAY(0 to 15, 0 to 99) OF std_logic; 
  											 
 
 
CONSTANT char_L1 : Screen_Line1 :=( 
 --///////////////Line 1/////////////////////////////////////////
('0','1','1','1','1','1','1','1','1','1','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','1','1','1','1','1','1','1','1','0','0',
 '0','1','1','1','1','1','0','0','0','0','0','0',
 '0','0','0','0','0','1','1','0','0','0','0','0',
 '0','0','0','0','0','0','0','0',

 '0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
--////////////////Line 2//////////////////////////////////////////// 
 ('1','0','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','1','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','1','0','0','0','0','0',
 '0','0','0','0','1','0','0','1','0','0','0','0',
 '0','0','0','0','0','0','0','0',

 '0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0',
 '0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), 
 --////////////////Line 3 ///////////////////////////////////////////////
 ('0','0','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','1','0','0','0','0',
 '0','0','0','1','0','0','0','0','1','0','0','0',
 '0','0','0','0','0','0','0','0',

 '0','0','0','0','0','0','1','0','0','0','0','1','0','0','0','0',
 '0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0'), 
 --////////////////Line 4////////////////////////////////////////////
 ('0','0','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','1','0','0','0',
 '0','0','1','0','0','0','0','0','0','1','0','0',
 '0','0','0','0','0','0','0','0',

 '0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0',
 '0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0'), 
 --////////////////Line 5/////////////////////////////////////////
 ('0','0','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','0','1','0','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',

 '0','1','0','0','0','0','1','0','0','0','0','1','0','0','0','0',
 '0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0'), 
--////////////////Line 6////////////////////////////////////////// 
 ('0','0','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','0','0','1','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',

 '0','1','0','0','0','0','1','0','0','0','0','1','0','0','0','0',
 '0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0'), 
 --///////////////Line 7//////////////////////////////////////////////
 ('0','0','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','0','0','1','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',

 '0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0',
 '0','0','0','0','0','0','0','1','0','0','0','0','0','1','0','0'),  
 --/////////////Line 8/////////////////////////////////////////////
 ('0','1','1','1','1','1','1','1','1','1','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','1','1','1','1','1','1','1','1','0','0',
 '0','0','1','0','0','0','0','0','0','0','1','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
  '0','1','1','1','1','1','1','0',

 '0','1','0','0','0','0','1','0','0','0','0','1','0','0','0','0',
 '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'), 
 --////////////////Line 9/////////////////////////////////////////
 ('0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','0','0','1','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','1','1','1','1','1','1','0',

 '0','1','0','0','0','0','1','0','0','0','0','1','0','0','0','0',
 '0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0'), 
--/////////////////Line 10/////////////////////////////////////// 
 ('0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','0','0','1','0',
 '0','1','1','1','1','1','1','1','1','1','1','0',
 '0','0','0','0','0','0','0','0',

 '0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0',
 '0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0'), 
 --//////////////////Line 11////////////////////////////////////////////
 ('0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','0','0','1','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',

 '0','1','0','0','0','0','1','0','0','0','0','1','0','0','0','0',
 '0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0'),  
 --//////////////////Line 12///////////////////////////////////////
 ('0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','0','1','0','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',
 
 '0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0'), 
 --///////////////////Line 13//////////////////////////////////////
 ('0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','0','1','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',
 
 '0','0','0','0','0','0','1','0','0','0','0','0','0','1','0','0',
 '0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0'), 
--////////////////////Line 14///////////////////////////////////// 
 ('0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','0','1','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',
 
 '0','0','0','0','0','0','1','0','0','0','0','0','0','1','0','0',
 '0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0'), 
 --////////////////////Line 15///////////////////////////////////////
 ('0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','0','0',
 '0','0','1','0','0','0','1','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',
 
 
 '0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0',
 '0','0','0','0','0','1','0','1','0','0','0','0','0','0','0','0'), 
 --/////////////////////Line 16////////////////////////////////////
 ('1','1','1','1','1','1','1','1','1','1','1','0',
 '0','0','1','1','1','1','1','1','1','1','0','0',
 '0','1','1','1','1','1','1','1','1','1','0','0',
 '0','1','1','1','1','1','0','0','0','0','0','0',
 '0','1','0','0','0','0','0','0','0','0','1','0',
 '0','0','0','0','0','0','0','0',
 
 '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
 '0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0')
 --/////////////////////////////////////////////////////////////////


 ); 
 
							 
variable Line:integer:=0; 
variable Pixel:integer:=0; 
 
	begin       --initial the screen 
		if Clk25'event and Clk25 = '1' then 
			if (Horizontal_Counter >= "0010010000" ) -- 144   why from 144? 
			and (Horizontal_Counter < "1100010000" ) -- 784   640+100 
			and (Vertical_Counter >= "0000100111" ) -- 39     why from 39? 
    		and (Vertical_Counter < "1000000111" ) -- 519     480+39 
			then 
				Red_out <= '0'; 
				Green_out <= '0'; 
				Blue_out <='0'; 
				-----Line 1	 
			  	-- if (Horizontal_Counter >=  "0110111000" )--440    640/2-24+144 
			  	if (Horizontal_Counter >=  "0110111000" )--440    640/2-24+144 x
				--  and (Horizontal_Counter <= "0111101000")--	488    640/2+24+144 
				and (Horizontal_Counter <= "1000011100")--	488    640/2+24+144 
				  and (Vertical_Counter >=	"0011101000") --232      240-8   y
				  and (Vertical_Counter <= "0011110111") then -- 247  240+8-1 
				  	if(Pixel <= 99) then --Line 1 Lets make our Text WHITE 
				  		 Red_out <= char_L1(Line, Pixel); 
						 Green_out <= char_L1(Line, Pixel); 
						 Blue_out <= char_L1(Line, Pixel); 
						 Pixel:= Pixel+1; 
				 	 elsif(Pixel >= 99) then  -- All else BLACK 
				  		Red_out <= '0'; 
						Green_out <= '0'; 
						Blue_out <= '0'; 
				  	end if; 
					end if; 
					end if; 
			if (Horizontal_Counter > "0000000000" ) 
      		and (Horizontal_Counter < "0001100001" ) -- 96+1   generate the hs_out and the vs_out 
    			then 
			  		hs_out <= '0'; 
    			else 
      	  		hs_out <= '1'; 
    		end if; 
			if (Vertical_Counter > "0000000000" ) 
      		and (Vertical_Counter < "0000000011" ) -- 2+1 
    			then 
      			vs_out <= '0'; 
    			else 
      			vs_out <= '1'; 
    		end if; 
 
			Horizontal_Counter <= Horizontal_Counter+"0000000001"; 
    		if (Horizontal_Counter="1100100000") then    --800? decide the frequency of Hs 50000000/2/800 = 31.25K Hz 
      		Vertical_Counter <= Vertical_Counter+"0000000001"; 
      		Horizontal_Counter <= "0000000000"; 
				Pixel:= 0; 
				if (Vertical_Counter >=	"0011101000") -- First Line  232 
				   and (Vertical_Counter <= "0011110111") then     --247   
						if (Line <= 31) then 
				  		Line:= Line+1; 
						elsif (Line >= 32) then 
				 		 Line:= 0; 
						end if; 
				 end if; 
    		end if; 
    		if (Vertical_Counter="1000001001") then		--521?  decide the frequency of Hs 50000000/2/800/521 = 59.98 Hz   
      		Vertical_Counter <= "0000000000"; 
				Line:= 0; 
    		end if; 
  		end if; 
	end process;	  

end Behavioral;

